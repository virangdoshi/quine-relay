module QR;initial begin $write("%s",("let s=(\"Module QR:Sub Main():Dim s,n,i,c As Object:n=Chr(10):For Each c in\\\"<?xml version='1.0'?><?xml-stylesheet type='text/xsl'href='QR.xslt'?><xsl:stylesheet version='1.0' xmlns:xsl='http://www.w3.org/1999/XSL/Transform'><xsl:output method='text'/><xsl:template match='/'><![CDATA[sub f(s$,n)print(s$);:for i=1to n print(\\\"\\\"\\\\\\\\\\\"\\\");:next:end sub:f(\\\"\\\"write,format=\\\\\\\"\\\"%s%s%s%s\\\\\\\"\\\",\\\\n(\\\\\\\"\\\"\\\"\\\",2):f(\\\"\\\"write{-}{txt}{echo -E $'(\\\"\\\",1):f(\\\"\\\"\\\\\\\"\\\"with Ada.Text_Io;procedure qr is begin Ada.Text_Io.Put(\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"trans B(Buffer)\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"trans O(n)\\\"\\\",2):f(\\\"\\\"{\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"B:add(Byte(+ 128 n))\\\"\\\",2):f(\\\"\\\"}\\\"\\\",9):"));
$write("%s",("f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"trans f(v n)\\\"\\\",2):f(\\\"\\\"{\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"O(+(/ n 64)107)\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"O(n:mod 64)\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"O v\\\"\\\",2):f(\\\"\\\"}\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"trans D(n)\\\"\\\",2):f(\\\"\\\"{if(< n 4)\\\"\\\",2):f(\\\"\\\"{f(+(* 6 n)9)48\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"{if(n:odd-p)\\\"\\\",2):f(\\\"\\\"{D(- n 3)\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"f 27 48\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"f 36 11\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"{D(/ n 2)\\\"\\\",9):f(\\\""));
$write("%s",("\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"f 21 48\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"f 48 20\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"trans S(Buffer\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"STRINGz:=REPR226+REPR153,a:=z+REPR166,b:=a+\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"2\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"+z+REPR160,c:=b+\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"8\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"+z+REPR165,t:=\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"class QR\\\"\\\",2):f(\\\"\\\"{public static void main(String[]a)\\\"\\\",2):f(\\\"\\\"{a=(\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"write(\\\""));
$write("%s",("\\\",4):f(\\\"\\\"'implement main0()=print(^1^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"BEGIN\\\"\\\",2):f(\\\"\\\"{print(^3^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"echo ^1^\\\"\\\",4):f(\\\"\\\"'f(s)\\\"\\\",2):f(\\\"\\\"{System.out.print(s);\\\"\\\",2):f(\\\"\\\"}s=^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"389**6+44*6+00p45*,^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\";for(c:(^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"#include<stdio.h>^8^nchar*p=(^15^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"Ra#include<iostream>^16^nint main()\\\"\\\",2):f(\\\"\\\"{std::c"));
$write("%s",("out<<(^31^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"class Program\\\"\\\",2):f(\\\"\\\"{public static void M83abbSystem.Console.Write(^63^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"Quine Relay Coffee.^64^n^64^nIngredients.^64^n^63^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\");for(int i=9;i++<126;)[3pva$^63^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",2):f(\\\"\\\"{i\\\"\\\",2):f(\\\"\\\"} g caffeine \\\"\\\",2):f(\\\"\\\"{i\\\"\\\",2):f(\\\"\\\"}I3b54rja^64^nMethodv4f#aeach(char c in(^63^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\")))^127^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\"));
$write("%s",("\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\")^127^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^32^[2al3dp3c[2cs3c,3l[2k@3kqa^31^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\")s rts(ecalper.h3eja^127^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"     53c4a SUTATS(egassem^127^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"rts(nltnirp(])]^127^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\".NUR POTSu4cba.C3dh3dX3bba[65bX4df5lga\\\"\\\",2):f(\\\"\\\"};)06xm3f$3loa)1(f\\\"\\\",2):f(\\\"\\\"{#qp]^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\""));
$write("%s",(",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'[p]#3sv3r23)ga3(f\\\"\\\",2):f(\\\"\\\"{#.33)ba7g4-ba5R4w23F&7d33&q7u53sda,4353.ma^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"' D ; EYB RCL4/v4+ja13(f\\\"\\\",2):f(\\\"\\\"{#DNEm4[m4ada. A~5[p4deaPOTSn4[#5e~5[o4boaRQ margorp dnex4[x4abaS*5[m4c2<[ba9i4[i4dba&#6[k4agaS POOL&<[77dba^1"));
$write("%s",("^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'j4[j4[j4gda&,)(6[<>cga. TNUO<7[s4bfa(rahcf:[(5dgaB OD 0?>[t4cca&,+<[ha9(f\\\"\\\",2):f(\\\"\\\"{#)A26[9=d4=[,6cqaEUNITNOC      01z4[a9c,5[U8dJ7[WFeeaRC .p4[p4aka,1=I 01 ODt4[OKecaPUq4[*I[5<gva;TIUQ;)s(maertSesolC;dYe$4Rra322(f\\\"\\\",2):f(\\\"\\\"{#tiuqn\\\"\\\",2):f(\\\"\\\"})652=5[qa^32^\\\"\\\",2):f(\\\"\\\"})974(f\\\"\\\",2):f(\\\"\\\"{#n\\\"\\\",2):f(\\\"\\\"})215iY3b8,ya99(f\\\"\\\",2):f(\\\"\\\"{#etalpmetdne.n\\\"\\\",2):f(\\\"\\\"})4208[.zX3ca02-Y[v3bda116~K[-L[j4ldamif+6[ga)30341\\\"\\\",2):f(\\\"\\\"}5[,6[j4lbat(6[(6c%a315133A71/129@31916G21661421553/04[04c(a%%%%\\\"\\\",2):f(\\\"\\\"}*+1%%%%811 -\\\"\\\",2):"));
$write("%s",("f(\\\"\\\"})48361(f\\\"\\\",2):f(\\\"\\\"{#j:+1 j@34[34cbawm4[m4cl4[l4cbaWm4[m4cba\\\"\\\",2):f(\\\"\\\"{m4[m4cva)(esolc.z;)][etyb sa)t=[#>[j4[~Jjca69m4[x5[j4lba,l4[w5[j4hla!\\\"\\\",2):f(\\\"\\\"})23(f\\\"\\\",2):f(\\\"\\\"{#~~v4[%5[j4hea(rt.o4[z5[j4hba)A7dda\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"};l3efa~~dneo3hra~~~~PUEVIGESAELPnr3ala~~1,TUODAERw3a63j$a(etirw;\\\"\\\",2):f(\\\"\\\"};u=:c;))652%%%%)u-c((||13jda#-<q3jda||i)3mhaBUS1,ODs4qka)3/4%%%%i(N4cx5kU4xPa2=:/t;2%%%%t+2*u=:u\\\"\\\",2):f(\\\"\\\"{od7 ot0 yreve;i-=:u;1=:+i\\\"\\\",2):f(\\\"\\\"{od))1(evom(dro=:t elihw?s;)s*45oi5vv3jd7dladohtem dne.s3dganrutern3d~aV);gnirtS/gnal/avajL(nltnirp/+Za|atnirP/oi/avaj lautrivekovniJ3d.4j[2cib\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"};0=q;)]q[c=z(tnirp.tuo.metsyS;)0(tArahc.y+z=]++n[c;y:]q[c?n<q=y\\\"\\\",2):f(\\\"\\\"{)"));
$write("%s",("0>2%%%%++i(fi;48%%%%)31-)i>3c&as(+87*q=q\\\"\\\",2):f(\\\"\\\"{);81312<i;(rof;n)rahc(+K4r[2k*3&oa=]n[c);621<n++r4aqa0=q,0=n,0=i tni;N3&oc6agi4asdRbQeclxfvfVk?f<bedRbzkF-;agb-a|dzdxd?fGb8aqeRdYd5a\\\"\\\",2):f(\\\"\\\"{b2b5i;agb-epb>aqeRdHa>aJaRaAdteFbae:b6aOa5aac1g\\\"\\\",2):f(\\\"\\\"{fyb9aS*4aLa7a;a4a<a=hcmkdxd;aNa?c6a|eebHaFaIaebzeJaeb9a/a6a2dQbUe-f2a-f9aS*5d6cRbC3gUc-f/aof0f?fSg7e\\\"\\\",2):f(\\\"\\\"}h4e.b2e6aRa;d2MVf4A5h;aTapc4aLcEegiof6amc6a-f;f:lsbdh/RDfybxcxc>aGaUeAa2a6ajg7a6a@ahg:a?aMbKaKa6a?e:a362aigGfMbIfTh>a:b1angamBf\\\"\\\",2):f(\\\"\\\"{bHa4atc3is5rjC-wbEc51JaMa\\\"\\\",2):f(\\\"\\\"}bJaDYEc-bJaJaUa-bJaMdJa8b7,;a1wTaKa1wTaP\\\"\\\",2):f(\\\"\\\"}rj\\\"\\\",2):f(\\\"\\\"}bE2W2NawwKa1wE|Ta1w1wwGs5wb\\\"\\\",2):f(\\\"\\\"}bJaLaJa8bq6s5h4c\\\"\\\",2):f(\\\"\\\"{a8bs54bs5:b+bC-rjC-rj\\\"\\\",2):f(\\\"\\\"}bJaHa\\\"\\\",2):f(\\\"\\\"{3a;"));
$write("%s",("3a-aHaJaFdQy;a8bIt:aUa:a7,di@f>fBl4ay6sbsb2be3^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'madiDa-a|bW*-a>6aua?aGaUe>avjhgKaKaigGf~6cgaHf?jRf&6esasbdh*b-a/bxcHa|f>ke3c2c\\\"\\\",2):f(\\\"\\\"}bhgXghgcg1ang\\\"\\\",2):f(\\\"\\\"{bHa>k?f-e:a:a\\\"\\\",2):f(\\\"\\\"}bHa?ahgJa\\\"\\\",2):f(\\\"\\\"}b5aAdte@a1angri>kxcpb7anb2b:bhg2f.j@dCf6aNjxcHaSfQfOfVj-aBfrifi?f-fng@f|f>kzeAgfiHaLj;a/a2h<bmhEh<apb/a2hEhnb<a\\\"\\\",2):f(\\\"\\\"}q:bhg/awh:fnglgFani|b1aTh3b:bhgJa7bHa>kHaUeoiCe|bxc3b0a:bhgIa|bzeJa|e5buaQbfi<b=a-a9m*c3bxdUem3aea|b9ai3eta2bMa7aZg|bXgVgTgRg9m3bIauTSgKcdc/bPcgfvf<h:X7aEa|b*k|kMa9m*cEc,dJa>a2a:b6agjykMa9m|b*i+cJ"));
$write("%s",("h6a33ifb|b*ir+|Jyg/a2h=aXhRalbOaCdlbOakbUagbRwXh1kDh7b5aLj?fwbjjUe2b5azgFi4b-bhcUrRjRjEu0c/bxd+h\\\"\\\",2):f(\\\"\\\"}hVi7?aea6a2bZ>ewc|F+F6azn2a5a*lrNjg3hQk?9xjDhBhgnHa1dmd9h?f1k;kHa:e1k;k+l<b3bxd6a*h5k=hmdHRShShxb\\\"\\\",2):f(\\\"\\\"{iacPa;a,b<hdufbpbubldic+d,bnbWfbjZiQh7-\\\"\\\",2):f(\\\"\\\"{jGkchEkuj<b<b<b4j:b*j<b<b,c9j6j7b-b9jXNAg3bDduk;i9a7bwg-a5bP|,c9j=a9a7bubxbs3e33eca1j33eea.bxkE3c33igaJb7bKf^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'3eka1jXNEj9a8*)3aoa.bIXjkWi4k,c9ji3a=aZlPg.bNg,c9jsb?fTjPk:k:i2jCa:i6aTjPkQjuj6aHk0kHjOksk<bze[CceaHajgS5cca,k53cGa:k8k3a6a<bShJiqN2b2a2anLNjJkriwbjj?f6Inc:"));
$write("%s",("e7b5aDf=anbNjybnk5a,bJa6aqAa^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'aubJa7b5aCgwbjjHa:e-b9a9b9aYjNjfg>am3awa@a@aNjfg6I:a|b9a0b9a6IVBamb>e|b>g9bJa0bNjfg-b9aYj9aCaAaJa9bNjnbJa6a|b5a,b?f:e-b*k-<-aRg9apbEuw3aRdinLfg8bAd5h-anL*b.bbb-anLfg7u3j5anLKc,i8Nxd6a-b9a8b9a7bJcJaybzm>aSh>aJa*c@dxc?b?so3a3a-b9lteUe6I<a2b5aDcxbvb:atcJaub5aEcxb7-,b4b-bDgi;aiaDkBkmd9h-7goaNkLkpb;awbjjnlo5a<bw3*D:Y|D8YJdHdplwn:n3lWl*n|nunn--n.bN8bT7K/xN44w=Q+|XwjbFnKxjkDYrst=jb*I.b<FvbEWI<0vZaZn\\\"\\\",2):f(\\\"\\\"}Plbo6ZaZn*oy6,bLqkxOoSaZuz21b?+>a\\\"\\\",2):f(\\\"\\\"}p?egB>a@X;Mg3ibKnD\\\"\\\",2):f(\\\"\\\"}84c*dAaYa/@ETAaUujbDai"));
$write("%s",("w?+@Xjb\\\"\\\",2):f(\\\"\\\"}=DaibPa*\\\"\\\",2):f(\\\"\\\"}fXxbZskbRzhXu6G.\\\"\\\",2):f(\\\"\\\"}y6QEa1bu9W9lbw>+1=aXa9v3b=|ioEakENto0TDAaBa3/vbl-I<<|3ob@ptctC|Za-b5|jkguWart*\\\"\\\",2):f(\\\"\\\"{L\\\"\\\",2):f(\\\"\\\"}qwwgA\\\"\\\",2):f(\\\"\\\"{Q+,o*x-b<ResPa>a@RA1XV9DfbgMd|zb9Dvbp2ossg1zHR1F+C3N9b3b*bhb;+kbRBWEfN6btK8zU1r0bTo5gbjbtbg\\\"\\\",2):f(\\\"\\\"}YJazS2Ir::/uOHwbN>W52pn5J7|9-R61hqXa-2,3jkFa*QL\\\"\\\",2):f(\\\"\\\"}EabPNa3:|rRAnYQ5kb:.26e.dI*KnSaEwN/PrTKTarr|oysYn;:jb1\\\"\\\",2):f(\\\"\\\"}8bvyC=Ua;:T.nT4bFa@yQE945iLsL|f7B,L:=anA3>CuEop\\\"\\\",2):f(\\\"\\\"}XnNv\\\"\\\",2):f(\\\"\\\"{ysqSaH;Gag.jbh4Kq>a-:-yTxjbgBjb4bxunvjb0b|\\\"\\\",2):f(\\\"\\\"}CaM=3bxxdb3jzAV*Va1/H,T|STcbwMShh=CSxv*-lb5b.bH,d*kbs5YnDncvG.P*Wn97EaLH,bST<a,b8b5b6b91zAAaYa/*0bOaR-AalRE?=s<rEadbwbwr\\\"\\\",2):f(\\\"\\\"}0hoc+NtA2>a>r*btR\\\"\\\",2):f(\\\"\\\"{bhB>rz7,3a7\\\"\\\",2)"));
$write("%s",(":f(\\\"\\\"{b1Pjblt@atqjbC0YR=p;pmbbP66e3a:\\\"\\\",2):f(\\\"\\\"}YaI\\\"\\\",2):f(\\\"\\\"}Da>aaKo2HE*bTag>93;o@pvbu|+wQ;uuSu>a1.b6#3aUciw*b5ACRkbfhP*6Y932pjbZa=OI\\\"\\\",2):f(\\\"\\\"{DaRAbu1;X\\\"\\\",2):f(\\\"\\\"{jbDaAaUJmblbDavbs8CIK?VYb@\\\"\\\",2):f(\\\"\\\"}iUnIKlbBaDnb+EawbDaux9bKpvp<aE9IS5C9bKpfOv2kbSa+,a-jbShYNv2ss,baznDao2bsrONaou-iwzbXnmbwTSh;LSajbDYS,;oIrazhbTatPhqjvTnyoH|V>Tn6bb+Ea0AfN?OTaDwZafX.PTn8blbBaEa6b\\\"\\\",2):f(\\\"\\\"}vazP|aoC0\\\"\\\",2):f(\\\"\\\"}rP|azaJGNFn0pSajb:6e?cFa30d<\\\"\\\",2):f(\\\"\\\"}UBaEa|bECWXo6DwoRvp<a2pB,=aE9=qC,d08o.bFnvpDaTa\\\"\\\",2):f(\\\"\\\"}rFnvpBq\\\"\\\",2):f(\\\"\\\"}ormB,,;gb-@1baK|:pWhb1bgbjb6b;p<r2My\\\"\\\",2):f(\\\"\\\"{u\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"{sDaVVyC0X8|02|M=a8oQptbwMOXtMmI*b,vjM\\\"\\\",2):f(\\\"\\\"{rP*?el0?\\\"\\\",2):f(\\\"\\\"{vbfR6p7b=a*bjM@aLraMVpk<;|,6Vp>+mIT<,bV3Vaec=p\\\"\\\",2):f(\\"));
$write("%s",("\"\\\"{b/P>Y<qVa4bY:cvUpr-J>=aTa<qNaVg9y<*#3a9aecSDu*1;*qQpp\\\"\\\",2):f(\\\"\\\"}VXTa4A<J0b1;7,RnDsrETaI5z>CBQImGRPib8**6e=ahukbhBjb:7Za2<hbqpYMBaizGhKKIKDaGKabEKUTCK,i@KDaCK8b4bCN33a2by78K6K:7kVt4EP+o/oF8abouB>|Xmy<a?ei9q0CsN4@yD,RaE*>a5potc.Z-S\\\"\\\",2):f(\\\"\\\"{OaDsab=atR+bj<<qZ*s5j<<qlb*pE*>a7rebBaKq=axuMkTaGNIEryP4hbVaD=28YaVaDE$4adb1bK\\\"\\\",2):f(\\\"\\\"}1bFay6vQ3EO+yb\\\"\\\",2):f(\\\"\\\"}<TsabOaC8l<+7Kty6ebXaWvvQy6jb1bXP@aGN2bZaDtFa@wU9Y*j63Aj6PB<jgH:.p\\\"\\\",2):f(\\\"\\\"}3b=X*6eudZ*|@zb\\\"\\\",2):f(\\\"\\\"}b\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"{DyEpK>IW7pWxh\\\"\\\",2):f(\\\"\\\"}Sh8Byxuv*b-+ldZA4b*bYs;ywoIyShvqZsQ<gtGaHXF4Zafb28qoW5g3Aa+,O17mN\\\"\\\",2):f(\\\"\\\"{i90b-<zWd2:g<xJ;Nw?2OaYUVDTKwrHWYab;fCmviq\\\"\\\",2):f(\\\"\\\"}MbOes6b5b\\\"\\\",2):f(\\\"\\\"{*7A73|<Xa;5hPBaNQKx\\\"\\\",2):f(\\\"\\\"{N\\\"\\\",2):f(\\\"\\\"}9sgOqSa>rO"));
$write("%s",("7BSGwPwU2LH,YLQ=0iwZ*qT6r/U2pxw\\\"\\\",2):f(\\\"\\\"}<GaeAq*DxH,v9bEzbdb6zSh>qzbO+iqGa.XtrsyjbH/2Bcvi9?w2pjd=a\\\"\\\",2):f(\\\"\\\"}b?aOEYRc\\\"\\\",2):f(\\\"\\\"{fbk\\\"\\\",2):f(\\\"\\\"}j7vu=fvd,bL,LAz=11j+s5*be\\\"\\\",2):f(\\\"\\\"{2rUaI<EC/U5bjLe|u<cbeBBajBr-r::gH+os\\\"\\\",2):f(\\\"\\\"{bwsjbft\\\"\\\",2):f(\\\"\\\"}/Yf,b07.7IXpYYaJ4YFc5KG2;+bO<U\\\"\\\",2):f(\\\"\\\"}wbJzdsy6M0Y*.KM0AqFn>r9b0ZFa7.IqT|R|*b1NL:RPzbbby74b4wTa1zn8Za7FMtV/tbzbGz2pzEV7Va+??A2pN;fLJpOV<\\\"\\\",2):f(\\\"\\\"{o@@<VQ2vhb@vShetkbebZa@Mp.9b8r70BaGCQ<+yN;Wq/B-bSqK>Oz|omxZ7zEV7AqMfsr|bQ>iF9<Gak4jby;@auh~6e0bS62vzbU4?ZebxxSaAz=aSc>aWnwZdb2\\\"\\\",2):f(\\\"\\\"}lzmRM.Da|Tjd>WE*-<fR.s\\\"\\\",2):f(\\\"\\\"}|U31*xbZa1bC|i48Acqubnu.s\\\"\\\",2):f(\\\"\\\"}|qU/7ib;|Vf1bT*6bibivT5C|Nk**2|NXIrxRS<ttcAs5L;au%3e=aS<ttb+Ga6=DOT*dbL*3bDO/72k*LTm\\\"\\\",2):f(\\\"\\\"}x@tzO?rE:@/3u8|dbHp"));
$write("%s",("K52bv,w3aWa+T80dbbbYfI:=\\\"\\\",2):f(\\\"\\\"\\\\\\\"\\\"),\\\\n(\\\\\\\"\\\"{rhAaShK*fh8AZa-bGazCf>\\\"\\\",2):f(\\\"\\\"}9psOrz8\\\"\\\",2):f(\\\"\\\"}9.4=AP*xRrtpt5V|q5|8bXaW-OiZ1PaztUadt$6e/ajbIVebiv-bSarjDaOa7*@=.K9bCa3KL7-dqvKqJ>wrI3aMc3sQ>eC:za=Q>eCFR0\\\"\\\",2):f(\\\"\\\"{Ta6bV\\\"\\\",2):f(\\\"\\\"{>=?aJ;Z.zw4/ct*r7.ybV\\\"\\\",2):f(\\\"\\\"{I/wbQIiwibCxV\\\"\\\",2):f(\\\"\\\"{I/huBt95.r4wC+ADkb2Mct2bbbCamzgMM0nKFRsp*p-bn-g>8miwib0bAtkXGzb,Z+AvPaGw<aWa*b.brZEwC+4\\\"\\\",2):f(\\\"\\\"{Oaj38C-EAa|*tY+\\\"\\\",2):f(\\\"\\\"{NaEaQ7Ar>8zb2blbU.1b0v8bkwTa\\\"\\\",2):f(\\\"\\\"{-cby-cxqZUagb@6|.qZVC+oo:<LqLmps\\\"\\\",2):f(\\\"\\\"{f:6byKzd9r3jnKJznK<x.6epd\\\"\\\",2):f(\\\"\\\"}NxuXwLW?J.dE|\\\"\\\",2):f(\\\"\\\"{w+b|.8v1bxt\\\"\\\",2):f(\\\"\\\"{bqYOJBLPWSqFsoRiblj6?YaLq90.r3ozsV.d2DtEawb<ad<6qdDSaldQaP<+?kbjFx2jb0bNF<aOaGaZqXqzLICmMIhcbB1QFTa/bb>C+fIq-/pybcb:ThqfIu0j1UqX"));
$write("%s",("a4TMo|b0\\\"\\\",2):f(\\\"\\\"{qoU7CalIP=dbjb.uUy1bwbgv*\\\"\\\",2):f(\\\"\\\"{v1E2JLC1mR=s+7S;2b+\\\"\\\",2):f(\\\"\\\"{N0E;b@3r6b-9s\\\"\\\",2):f(\\\"\\\"{m1\\\"\\\",2):f(\\\"\\\"{b,Pe>s\\\"\\\",2):f(\\\"\\\"{g9kbk0t0,dJ-T\\\"\\\",2):f(\\\"\\\"{E?,3xbssRn\\\"\\\",2):f(\\\"\\\"{OCn>=8bowb\\\"\\\",2):f(\\\"\\\"}>Hq-4Ox6eSaXs-Yg=sr@aGqitdERXhDjb*-@XRao63s9/0FD|8bvF73hBYuTao6Oa\\\"\\\",2):f(\\\"\\\"}L|S9rp=hbn*F|9/wbDysh4b13cxbBw3K3vbO6|;<72cbVa3ba6T|YFr6d:Xshxhb7b2.mo/b+s/y0z=-wrjjoz*bB<Zaj-mbShx*s>q>Oia|gbcLVUJAZaETc9P/@-*b=-E;iqVV<|\\\"\\\",2):f(\\\"\\\"}Ka^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'aJrQvgkzofb0b<=Q5m3pTZ3p58bIoJAMvCvd4a6a9C+babhJGaw?+bUa11dK6bQan"));
$write("%s",("vJwr2ubNwJ48CBa6C*b80QaDE9fscY.E=ptntEar?K\\\"\\\",2):f(\\\"\\\"};xBSTsjbYaLSN|Ba9PVgGS3i9*yWdbPa9b2pHWYaC?K6EaQam2Xa8-vQzxST48n*\\\"\\\",2):f(\\\"\\\"}30bWEmbqYUq2qFoXa2pITabM>N4M>/bKxpz1?2bCaa2-hJ3@pGnmRxb7Z.b5ZQaQFpV<at/8*QaShetEYyb:1mOPwtY2F**Sa@Wx6h.;L<rtDz=bbYEalb\\\"\\\",2):f(\\\"\\\"}bNvs\\\"\\\",2):f(\\\"\\\"{9/0bR-QaW*-bMvb+ygDa*w=aeb-b1.2BlbxtrsGJ5;8=4/AaYSQa3bD=?zz<NaYFRaqEab+/ewCIYaI0lSOa3shsNaEa06e#albcb5ilukbGq+bRazdSh/yWn?397Va=3asa1bqtkbLv2puC0s\\\"\\\",2):f(\\\"\\\"{br2x4cBavx<xYa@abbo@G2stkbe?GC2pH?kbKrH1@XUnG?*btbC;N4Oa|bOaguNan-NaEA3bec-YAnl6?ytb+bmb@?2bf@6M61J7c;xb9b>adUebO+Wt\\\"\\\",2):f(\\\"\\\"}|I0eR-yRas\\\"\\\",2):f(\\\"\\\"{t7bb4A;oSabbgb3b\\\"\\\",2):f(\\\"\\\"{o\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"{S*lbtzLHbb5z=-GBP;\\\"\\\",2):f(\\\"\\\"}BQ,92PRmpwXUqDACSj6\\\"\\\",2):f(\\\"\\\"}>*p+d\\\"\\\",2):f(\\\"\\\"{bPa;yL*.1DA"));
$write("%s",("gk2qwb,=g=Fvt7=a7DisEvfJ\\\"\\\",2):f(\\\"\\\"}kJXY,<aIGybcvxbdblqzbOU:6cDbH,bwS8zwkbDqQsKnp+nvCaubFaX@UaGN2bAqkb5bL\\\"\\\",2):f(\\\"\\\"}U2?rS-l8>qcA?tB<db\\\"\\\",2):f(\\\"\\\"}subFa:7vGz8xx|r1tvD-biwQI8E;ueA=SFaRBkvTMTaPGQa?aO797wbp5kbWnzb;|LHn=xbDan5rt9A|r@?q|<ocro3a:b\\\"\\\",2):f(\\\"\\\"{b+uIWaJt+jb4byswbZukbECH+2bd|QaqIgvKz\\\"\\\",2):f(\\\"\\\"}subAucbsgsP\\\"\\\",2):f(\\\"\\\"{AzbzblA/2wsVa1b6-1MptU-?aWJl9\\\"\\\",2):f(\\\"\\\"}0Shh=Gow4Oau4qZPaRaBK<ayb3vVACvkbf>?ub+LWTzDYS,Oa\\\"\\\",2):f(\\\"\\\"{b2b2vv5n=SGfebSlSv5n=nq1bP\\\"\\\",2):f(\\\"\\\"{o5+bEaOw2pp57,*b<ah4n|P?8blAw*tbmyYyyyLvg@3b;BYaRyux:\\\"\\\",2):f(\\\"\\\"{K3Jz.s>qR=Hv*b?aUa:4n=stb4abaFb4b7bDa\\\"\\\",2):f(\\\"\\\"{b2t9tq*NaCRlSGqDa2bK5ZumbIQmIF@2b\\\"\\\",2):f(\\\"\\\"{b?aU@K+.;;JgzFR.y*,h7Vq2bV6d\\\"\\\",2):f(\\\"\\\"{zbuA*boGej>ae=@Rm=QIgbRa.2ubyb\\\"\\\",2):f(\\\"\\\"{bjbx<5t1snjU86bSa"));
$write("%s",("x<\\\"\\\",2):f(\\\"\\\"}9D\\\"\\\",2):f(\\\"\\\"{sAv<+b|vdyCP^127^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^32^[2fha\\\"\\\",2):f(\\\"\\\"})1(f\\\"\\\",2):f(\\\"\\\"{#v3mja51(f\\\"\\\",2):f(\\\"\\\"{#,4353(za199(f\\\"\\\",2):f(\\\"\\\"{#(ntnirpn\\\"\\\",2):f(\\\"\\\"})215(f\\\"\\\",2):f(\\\"\\\"{#)|4[|4aFa|blbuxccjbSh>qhbTadr6g;5\\\"\\\",2):f(\\\"\\\"{bk\\\"\\\",2):f(\\\"\\\"}B*ZajbOisrkb\\\"\\\",2):f(\\\"\\\"{bSNq4*w2b7A.dfhi9r<;5wbBr@f#a4w0w.w=awqVf1?6b+bYaYakbf>7ro6i3cIc7T\\\"\\\",2):f(\\\"\\\"{b2ber9,guyN+vDq+?3b++Kx2Blbx@.bPa/bmEiwQIO:<z=A97Do*b?af|,iQa|rrx@ZCqTDlAyb,r\\\"\\\",2):f(\\\"\\\"}AEU6bfbaAb,Zsf*CtpP<JjjZsf*6bD/RPzbnYSasYb\\\"\\\",2):f(\\\"\\\"}wb\\\"\\\",2):f(\\\"\\\"}?2pk-OaEw61uuy+qojbkxfxW*-bfzO;=H\\\"\\\",2):f(\\\"\\\"{bdb/b,vVaZado4iab6pL4EwPE:5i58y/b\\\"\\\",2):f(\\\"\\\"{wzb-osQ=N,bW:N425DM/5d:x5?av5o|@?PBjHevi7=txb*Q|6a*dLU"));
$write("%s",("l>w3aRj>Ya*Qe=X4W1QamQ?rGoF@2\\\"\\\",2):f(\\\"\\\"}vG2pCa\\\"\\\",2):f(\\\"\\\"{bRB7K<wwqvbBsGw0XGaZqkbO|ebZ|yt3bB/WaSal6Vah>O+qo:obb*wa7\\\"\\\",2):f(\\\"\\\"{b+dosWxVUnjz6H?u6F4Z>SaI:euC:h:hx?aejdl|bxqTK|*Czab3>OaxZ?rZn=G0,jbIYTKTazb9bzuzLCSub4\\\"\\\",2):f(\\\"\\\"{-<+bmRo|I59bRaBKA2;wYa\\\"\\\",2):f(\\\"\\\"}35K|MH8TK|*/RabJ\\\"\\\",2):f(\\\"\\\"}2saU,weuSTtEK4A,5bQatE0Sz8|*S*d<Dyxbkv1bYaR\\\"\\\",2):f(\\\"\\\"}DXB@ubuCDy4b=\\\"\\\",2):f(\\\"\\\"{C8<Pz9o7Gn<aeb70K9eXXi/a\\\"\\\",2):f(\\\"\\\"{fRqJ78bC6t:2/YUYX3:/br:B+jb\\\"\\\",2):f(\\\"\\\"}.:3zbg:e:i4<:M5a1czbg:=73A-M>t,*n*ys8:G:.ikbI/h:I:T|lvyUmz9AmzWgGC4|Tabwg:y6CaWa;?lvPxoiwbYa-wzbg:w:Ua\\\"\\\",2):f(\\\"\\\"}.5CM+F:4|ybYadq\\\"\\\",2):f(\\\"\\\"}Ih:I:y7I59AF:Aak.v2f6sqOamzGS1J?aUa5v+:=:-wNr\\\"\\\",2):f(\\\"\\\"}IzbPahx9Amz/Rl/?albmz*bTVUa@a+bwqI9Xsc6zbEnq-nKPajIVaWaSamoDaEa,bku1;+?|6e$dUajHa8Cxb"));
$write("%s",("TwrHWYaR5CSGL0bK4A,btQasgVaP?Mw*Qbb\\\"\\\",2):f(\\\"\\\"}=<L|qs;o6TDK=Vp:pffq0:h*JMrlScLmoPRCqs5rsmEfhc-\\\"\\\",2):f(\\\"\\\"{TmbTYa4cqm=Za-bSaY*kbN*NkjyghnBrsOa0=KO\\\"\\\",2):f(\\\"\\\"}+Au2LNanqUa13HRYaxbIhitybBaRajZ+CYa7bz=TKH8vbZ-?Kr--zd5bmbtfbjbO+Zai=i+*bS<ebpFP7>Egx1b,ODaEa8b|bdbwv3>mwab1b3P9bTKYsB,D|5Hz;bj0v-bBaSaIpoCVa@6H\\\"\\\",2):f(\\\"\\\"{Eaeb:3d6:3NaqE,6e~bcbRnwbYaUa.bQa@67br6=aP7:6a|8\\\"\\\",2):f(\\\"\\\"{O6BaSH3TIE.@U7q+fw:AJ;b+IW:vQaPaTaSh;F9Ds1Wps17b30>aJCH\\\"\\\",2):f(\\\"\\\"{8A+GSanBAaubDaTa6zh.\\\"\\\",2):f(\\\"\\\"}|9w?Z.yqzb4cubkbhr,bsz2pMfkb9\\\"\\\",2):f(\\\"\\\"}5riwvbyy2o1b\\\"\\\",2):f(\\\"\\\"{vI|OaiA5CJw1bwb0bb@DYMoCo\\\"\\\",2):f(\\\"\\\"{bd<,btr11N5@wkVyATaH17b*,yoH|B0ubw*owb\\\"\\\",2):f(\\\"\\\"}7bKzbb/xFa.@bZ4fAas5Ua2ONaTaSa2b/C:7tH|\\\"\\\",2):f(\\\"\\\"}3HRanU\\\"\\\",2):f(\\\"\\\"{uh0EzDsBsrwPrZu?3B/,,O;+dosbb7bP@"));
$write("%s",("iBbucWaP?Pt,68uwboz8wOt-:UZ.q:g6eUaL=J-yUo5+b++sr+b@vMvUnT\\\"\\\",2):f(\\\"\\\"{=-0q2t0tH3moNavbuh3*Yawq3b\\\"\\\",2):f(\\\"\\\"{b02LvmbWV@v3yV5YuAalS-Egu6b@aVqWTFaoR,k|S|+wbp5?avCRa\\\"\\\",2):f(\\\"\\\"}TlbZaWXct?ZO3a:bxbRMND4A6rdb7bYjxbgCK\\\"\\\",2):f(\\\"\\\"}UTsvB*Ea43<r2bt:EowbYaoiB,ICLvmbd9sQt52pbNsg=Zkb1bbM\\\"\\\",2):f(\\\"\\\"}s.s>qdQS*sq*bV>|bq0lSjb+b=aPawlX+:\\\"\\\",2):f(\\\"\\\"{iFP;DaPBN8+bEadz-gUE2p?a-Mdbu@VTdudvYawFmbfbejXn2bvbw0EcT/:\\\"\\\",2):f(\\\"\\\"{Tg2Lh.vq\\\"\\\",2):f(\\\"\\\"{bSX0AKD3b2v5ifN1Pbvld|vtrsyjb3bJ7wbBaEazc0CBaDy-+fIDacby6U4qr7bV8w.=E6bfbDa\\\"\\\",2):f(\\\"\\\"}bwb8|:6p?yq\\\"\\\",2):f(\\\"\\\"}X*TDs4eSa:\\\"\\\",2):f(\\\"\\\"{ID<|bbqrk\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"{8wDcK*oVaL3n//TAaBwk7tYcbAvz|Y=mpwXjbH;n;FaU\\\"\\\",2):f(\\\"\\\"{WanFD-p\\\"\\\",2):f(\\\"\\\"}Z+s4.xlbDtvQq6ho,9-:ioY:?8/XpSlv3*3JHBQI\\\"\\\",2):f(\\\"\\\"}wp"));
$write("%s",("v\\\"\\\",2):f(\\\"\\\"}wK>IW4CwbjbP+bc,bmx@aBumj/HjS-xk7i74Mb<|6c\\\"\\\",2):f(\\\"\\\"{au<Ggp1d<j-06kRP;=8yo:w:p9bu9aVcCa9rzcVa0BtE>rgkjoCzH8U7=aGL3o|ZybYa,p;J9E5@Oa-RNaDNb|rtnAlA9x1MXnPZ9xvbz7QaAa5bFRe,Kx;M3oE*IWsEvblb2blbj=-tWxgbvby7112ONaaxabr:6LXDor|@+b-9.d.G.d\\\"\\\",2):f(\\\"\\\"}tlbDLGUy\\\"\\\",2):f(\\\"\\\"}I\\\"\\\",2):f(\\\"\\\"}-v.|SaS\\\"\\\",2):f(\\\"\\\"}1bSa=7Cp-9R\\\"\\\",2):f(\\\"\\\"}3baba-dE@a|@wb0bioiK=aJdW:V5Sa=aEa-bwy\\\"\\\",2):f(\\\"\\\"{bhbwyt*wyn-cbfFXa>,o6fbOp:wQAosQAevLvaw=bpb|D8YfbP6p\\\"\\\",2):f(\\\"\\\"}P655QACa*Ior-r6LL7?9m5s8r:6L+YybF@5b.bsq@a/Lw>V56LZaG,Bagh2bDx5HDEeUhKV8mq@aq4Da\\\"\\\",2):f(\\\"\\\"}0Mw+b-bHH*hc3uLbQAecwLB>Mj5Ytb\\\"\\\",2):f(\\\"\\\"{A-b,bvbUavfS>fhnYTKE*9UvgCA;OUTUtibFaIWo50Z\\\"\\\",2):f(\\\"\\\"{b:TOa5b6bPag8Oa<0Fq/b=rkbsO7.-t3/fh7.qFlbd5fbvkhb0DT7X@IqLfzqPEg=|oe7mE?w*h*IV6FajvQZ3/TJibY\\\""));
$write("%s",("\\\",2):f(\\\"\\\"}qKxb3v:@iY2zFPaQEOE\\\"\\\",2):f(\\\"\\\"{bMEF4xbvb6o|b4bd73yFq@<pv2b2pqZPabb3b>aF0=akOEPsrrqtbYa1?qYjSQZp8ubU@\\\"\\\",2):f(\\\"\\\"}o7A3bDNENc--t0boG5bOJfx2\\\"\\\",2):f(\\\"\\\"}Pa/xUadr?wacjy-tB0RGVFvboRPaI|qVf@abOCtRs*e8z96fDaN;fbo|S|f:kZntGKNap*q1S*R|uZK+Jxlb+?\\\"\\\",2):f(\\\"\\\"}L6b2bz5Wamv.h<aQafbW9w;Bwdo?\\\"\\\",2):f(\\\"\\\"{|b48sPkw0bG,:1DYibBY?aKY6h98/bd<oyQ<<TM.YaXaTz9J.P5Awb|o1q-B<a,pjbRV0lS9Z;Q98Wp|1b>a:yY5j<rr.\\\"\\\",2):f(\\\"\\\"}|S5RVaCSPaIqLNZW9\\\"\\\",2):f(\\\"\\\"}5iLN8bsrBs1G2b\\\"\\\",2):f(\\\"\\\"}b/b2p*w5gkbL4Pa@,*ogbrt6VRavzR6=8kxwyWXRauC\\\"\\\",2):f(\\\"\\\"{b=aE/mbZaJ0,i4\\\"\\\",2):f(\\\"\\\"{Ca0b9,NpTK,bShwPgOcbgy>acb9bkV2bBwXaf<RaxbzbgbxbkH;\\\"\\\",2):f(\\\"\\\"{\\\"\\\",2):f(\\\"\\\"}x-9V/Y2<wxbSh085t6byqCanttby.?a0bLGJG-yA+0z.z,z+\\\"\\\",2):f(\\\"\\\"{Aa,Ny1Op6qTaZnxs9bV*EaN;8bY5N8>We@I\\\"\\\",2):f(\\\"\\\"}/"));
$write("%s",("GAti\\\"\\\",2):f(\\\"\\\"};yIo2/CSOCSV0bE<2s6bxbVsvbYa*7kTCaE?bt.bBTFagqfbgbD\\\"\\\",2):f(\\\"\\\"}-5MUZ0KUQae*mOgfXsH|I\\\"\\\",2):f(\\\"\\\"}r-dOjxZxE4C4xM\\\"\\\",2):f(\\\"\\\"}P4b.qp8gbZ3*7h<|v\\\"\\\",2):f(\\\"\\\"{fr+tA2<2b>HYu9U+SopIVyz\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}LVBV4|DOgQ2p?rArxu5b|bEacN8b-b8b\\\"\\\",2):f(\\\"\\\"{bJmCRxz:pGL;Ve|UalAMv5bE;:p<V:VAv+bg@>aTmD\\\"\\\",2):f(\\\"\\\"{\\\"\\\",2):f(\\\"\\\"{b5bi1Waqtot7R,,g@H\\\"\\\",2):f(\\\"\\\"{*+>xU-uh2i|Vc9@-04hxhsJFN\\\"\\\",2):f(\\\"\\\"{F+K+uby\\\"\\\",2):f(\\\"\\\"}+bguA-jb8b-h,MDsnuFa8*LrS,d8vvRIAQlb1znsL|NagbctzLMTpxfs=tt8h3D\\\"\\\",2):f(\\\"\\\"}*5\\\"\\\",2):f(\\\"\\\"}DD\\\"\\\",2):f(\\\"\\\"}SS-v2Ltolv*Q/boGyoxxysPAld02,r=\\\"\\\",2):f(\\\"\\\"{p\\\"\\\",2):f(\\\"\\\"{jwUaUnKxE|Br3o<qsjxwm<NrOs|Tc4AD:DlbhqLfVq+bVDgb:7K+NvL*CxUa|9aSXaS\\\"\\\",2):f(\\\"\\\"}1\\\"\\\",2):f(\\\"\\\"}RBT76D1A+rZaRa@afsybCaI5hKW3ib?@mb3/lbouYFp*"));
$write("%s",("I533<ojbqtBr7\\\"\\\",2):f(\\\"\\\"{5pLvdShbQ<<wbbtoV@CRCa+?L-U7Aah4|J/TL.bb-b5blvZx8C<asgzbv<xbab;o@ai=*h6pCsTaE|Ugbw/LCa,b.bp\\\"\\\",2):f(\\\"\\\"}|b2kxy9D4bL4xxEvE;LsTv<s,b:sZ-.b9bhbl\\\"\\\",2):f(\\\"\\\"{bRsJZQft4q>app8CkSSsz6v|6baK5bH<,Kq6Daxbt-;|Oa?aubZ|rPdrS>p\\\"\\\",2):f(\\\"\\\"{RK8w<,oz+qfhX-vbkbTm-qnKQaQEX4|bLnc\\\"\\\",2):f(\\\"\\\"{ibft:7>aDo*-GLwb81=af\\\"\\\",2):f(\\\"\\\"{RMdxXa\\\"\\\",2):f(\\\"\\\"}bhbEr\\\"\\\",2):f(\\\"\\\"}C-1CodyvbYsSa4biPOQAraq|\\\"\\\",2):f(\\\"\\\"}5.J4utTO?t.bU*1M*q\\\"\\\",2):f(\\\"\\\"}b2bxpoIjbhNFaYaX@hbzBRA0b2;sM2z/bO@m2do,IdbvDuqPBiR\\\"\\\",2):f(\\\"\\\"{Ngb|b*b1bdb6ueo,qJ73AZ3wFU*xbd1tthBOagbH7RAi+8bgpYa\\\"\\\",2):f(\\\"\\\"}b*|\\\"\\\",2):f(\\\"\\\"{Qnvgt:uab-bKrEuC.E7nPIr0beb=afsmq\\\"\\\",2):f(\\\"\\\"{bEpOEI<gP,\\\"\\\",2):f(\\\"\\\"{i9bbj6O:Ew5C81j-A1Yqy.yd\\\"\\\",2):f(\\\"\\\"{sN?+<LHhsAp|.\\\"\\\",2):f(\\\"\\\"}QpPfboGhbuCV8Xad"));
$write("%s",("stbBq=r=8iwt,Qajb3sPGPE.A3su/b?2pDq*NEok+9;BLkb@2ebM\\\"\\\",2):f(\\\"\\\"}EarvVsluPa6u@FguHtt-dbP\\\"\\\",2):f(\\\"\\\"}L\\\"\\\",2):f(\\\"\\\"}ebFs@t,2EJSI,bHpCaY:i+y65A0|t1\\\"\\\",2):f(\\\"\\\"}Nlz<r3H7bjbabY:y;F?R0D8>@t75s36qLL*Zacb,d.z3bIGDafJwbvbab*0?Nj<Ea.z;yJ*;yIqebxpwrBi\\\"\\\",2):f(\\\"\\\"}b,b4HgInLqNPap+J8OEbbH<Ux<qef>ahBabn5xzI0tqK4.bIGctZ?yxjM91N>C;3E=-SHn-h6h\\\"\\\",2):f(\\\"\\\"}i9g+v|>aKo13zt5N6bS\\\"\\\",2):f(\\\"\\\"{J83bnBybW?*b3bgBgz,\\\"\\\",2):f(\\\"\\\"}@aab<afbrmEaZaEaabdbNBC+FaWpXa8w|bfNqsfxUa3jI0U*OMgOQatpYa9,<=u/@=E<j6=\\\"\\\",2):f(\\\"\\\"{N8.b\\\"\\\",2):f(\\\"\\\"}N2pJK?aR6L;I0dzeb4/sr,bnD*?;EvbeF;o9wGamN\\\"\\\",2):f(\\\"\\\"}=p\\\"\\\",2):f(\\\"\\\"{lbsrADi=Q;Raw0kb+,grcK,b/bu+V>MLP.xp6bvbMLM>J*ejJ74bOawbaNEas1OaJ*4A,bZ0t@A.\\\"\\\",2):f(\\\"\\\"}FnLebDo+sr>NaJ*Cq1tUaGtfblt5AY*Mn6*lp5bcq:u3vj+ubGaS=\\\"\\\",2):f(\\\"\\\"}k<=fbrv"));
$write("%s",("5y@7cl|uGAis618bcbZa+blAzJFay;W=5,V3?axtCq1ABo<ahb\\\"\\\",2):f(\\\"\\\"}bYfxblbQt9*-hTa*-Vq02eb+b3bVqa3i1yb0bk\\\"\\\",2):f(\\\"\\\"}GFubAaGFY\\\"\\\",2):f(\\\"\\\"}S\\\"\\\",2):f(\\\"\\\"}4?DaVaUxhb\\\"\\\",2):f(\\\"\\\"}+<*/bCa<aF4Lr+bWad|buSaebE5tb?+mzTm5bzL4we.lbxB,b2bzLp?ebuba3osI/ub\\\"\\\",2):f(\\\"\\\"}oQaR|9yY,2pkbD98b4?\\\"\\\",2):f(\\\"\\\"}0Ba@ahb2bdb<aa3Xa?uef|1G:ib?a5okxwbP1Z|Jwbdq0u16?Lnq6nLIbqJ-b37dly\\\"\\\",2):f(\\\"\\\"}qE9bZ*rsQ2t,tbPvmI/xjbT*hBlIQa,b6bZavw?a>K-dX|hqPBEambR7FavKE5F5,b3bbm.q\\\"\\\",2):f(\\\"\\\"}bybNpVfY=<5w\\\"\\\",2):f(\\\"\\\"{Tp1b=adbXadb2/Tqq6?a\\\"\\\",2):f(\\\"\\\"}bAD6fvb8q7,wbkqiq3b=rpzVauuDaa3RJ7.cboy2b0Du*I*Y4\\\"\\\",2):f(\\\"\\\"}03/Bp5t:\\\"\\\",2):f(\\\"\\\"}<aab./Pait6b,y|b\\\"\\\",2):f(\\\"\\\"}0Da8bC;v<sg6bBaY5d\\\"\\\",2):f(\\\"\\\"}9E@wCuksSg3bJ4D9/qUE=zYaE3Cak.E*jb-bQ7u*Czub9vqm2b|b+7;-=o;o9oq\\\"\\\",2):f(\\\"\\\"}VaE4kws"));
$write("%s",("5vb2o9bn+w09A8oD\\\"\\\",2):f(\\\"\\\"}F7s@W0yHzb5bpB8/WaFa<||bfodo0bboLoBuackb-t+yOn\\\"\\\",2):f(\\\"\\\"{,:ggbs6JIlb?a8unuOsgr3ECn@<T7ybkqE=c\\\"\\\",2):f(\\\"\\\"{<|wbp9DpN7,+T7RDcH<|::o7g8@a>aU-e73gDF78SGh\\\"\\\",2):f(\\\"\\\"}mj>a*bcblbEa+b/>*-:oro4\\\"\\\",2):f(\\\"\\\"{4bfbJ82qW-BzQa1bCaDahbq4mbvGWt9-mbu*P|?aWq91-pjy/>7bcbro0>Vau9F@aEXaUappdbo2wbvzcbRvfFR|ju>aw*b:zA\\\"\\\",2):f(\\\"\\\"{bEafbJyNqh<jxs847,bSaGad3.@d|>,Ba7uH/so=-G4xrD4:*|lwHVo\\\"\\\",2):f(\\\"\\\"{FB468BaRnK\\\"\\\",2):f(\\\"\\\"}OibtX2Y\\\"\\\",2):f(\\\"\\\"}C-ejJAq-lB8|tbJ?A\\\"\\\",2):f(\\\"\\\"{\\\"\\\",2):f(\\\"\\\"}x0qo5N@5t4umzH1r-3gh\\\"\\\",2):f(\\\"\\\"}>3\\\"\\\",2):f(\\\"\\\"{bn5tbeB3itzlpybhuzb35QAI8iqGxhb-b3*W4@ant\\\"\\\",2):f(\\\"\\\"{bwb\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"{6<d*Pj?*Qn0Eo*X4I|tb:7?aRaS*@aQayo9b2zP5c5qoTB8bhbs|g81\\\"\\\",2):f(\\\"\\\"{*--b2kfbg=|bB6k+Rav6K/\\\"\\\",2):f(\\\"\\\"{b"));
$write("%s",("ADO=fbTaHxpF:/Uag-1be\\\"\\\",2):f(\\\"\\\"{1\\\"\\\",2):f(\\\"\\\"{A9lqosubAFRatb9/Mqm*H+b?7t=aPDqrnuq\\\"\\\",2):f(\\\"\\\"}Ea=a.bpv5vE52p6b*>hkI\\\"\\\",2):f(\\\"\\\"}or<aXsebxvEa*bVaTwibZ0a<n>Mu\\\"\\\",2):f(\\\"\\\"{D0lyD6b48hE\\\"\\\",2):f(\\\"\\\"{b,bwbdy?rq1hbmb+z-9ux0vp*Xa-bt:\\\"\\\",2):f(\\\"\\\"}BwbP*O7FrJ;+7p=::Gal+ew2pv+Hn+bNaab6b0/A3Bw.0<aTajbdtMq?atbhoizVs@/i/6byb8bkbS.mbP;k*q6xB=Cubb?>=mb;wd17b\\\"\\\",2):f(\\\"\\\"{pK5-+a83pJ9cu2\\\"\\\",2):f(\\\"\\\"{4\\\"\\\",2):f(\\\"\\\"{4s9\\\"\\\",2):f(\\\"\\\"}dr.bz,=amb5bC>Na-bF<p24oSt-zxy?a3tebOATa\\\"\\\",2):f(\\\"\\\"{bRAK>.bxyxbI|hbRafbqmlb7t>aw0.29v/.Eyf\\\"\\\",2):f(\\\"\\\"{PB7\\\"\\\",2):f(\\\"\\\"{;oP?gqsjNaV|1yeo@a8/S<tDDaZ>ebFrS;z7G6Vs|BSa56o/@Cq|l\\\"\\\",2):f(\\\"\\\"{s3R90lP9-luBWappZaYf6bICh<1r8\\\"\\\",2):f(\\\"\\\"{zbAa?\\\"\\\",2):f(\\\"\\\"{OaKrebpz?a=BBuurWaj7+bbvxy/bEylvDs>6P\\\"\\\",2):f(\\\"\\\"{2kWaq|\\\\\\\"\\\"),\\\\n(\\"));
$write("%s",("\\\\\"\\\"xqSa2\\\"\\\",2):f(\\\"\\\"}r|Cv|-Dalb:\\\"\\\",2):f(\\\"\\\"{.bUsUa*b;15q48rxp**:5*xb93ajvb-bUxCaNac|Wg>ru<.bFa@zho:tBa:|N*ybXkEsCsAs4s2bNaluZ.Yh\\\"\\\",2):f(\\\"\\\"{bzoQaL-?3E52/LoL<Oa1bAawbHB;o?ai+\\\"\\\",2):f(\\\"\\\"{yd<7tho<ambTaLf.bP7ebfbEaN>L+b,>BP;5bFaMoQzOahbWqFnos=0qz/bFacbRa2p<aVs-uVaHAwA<ac*9b9b?aVa\\\"\\\",2):f(\\\"\\\"{b9bL1lb\\\"\\\",2):f(\\\"\\\"}b1rRap*n*TaZ0sBO9q@OaLq4\\\"\\\",2):f(\\\"\\\"{P7+bMrAaH>1bdt>aDaEvwb*rjqs8Rwebd*8uL37bTv<<vbzbSaFal|ho9Y2qwbYqWauhl|,bL:UjNa01R<wrb|2ph4ybk6<+2\\\"\\\",2):f(\\\"\\\"}Oa/bzb>aPa1bRah0vb*bMnibyw,3JsQ/K,U6db+bhbF=\\\"\\\",2):f(\\\"\\\"{baw?|3bBa4w=axz0?hbhbubU*XnRadbh\\\"\\\",2):f(\\\"\\\"}56Ww<a?ao|uh|9M?zbU2CpVn0*ff\\\"\\\",2):f(\\\"\\\"{delQaz=tbkbu+i:G6jk4qN8Qa\\\"\\\",2):f(\\\"\\\"{sd|b|AaxbD84bB8-\\\"\\\",2):f(\\\"\\\"}8vxb069q7;K/5pabY\\\"\\\",2):f(\\\"\\\"}6>fb4>|qeb,b7bS2LwM+u*zbOi<+E<UaF0u+"));
$write("%s",("D\\\"\\\",2):f(\\\"\\\"}C7m>D7k>\\\"\\\",2):f(\\\"\\\"}b.b?rs**o-,I5/uEjfb4bEa\\\"\\\",2):f(\\\"\\\"{bS,0b.vFaR|7wqo.b7..>.utloz5bTmWawb|\\\"\\\",2):f(\\\"\\\"{Ta7bCqVa\\\"\\\",2):f(\\\"\\\"}bdbtbP<9b@/jqNaz=Ba,yZuWa6vf>it/3NaJ;gb/iY4\\\"\\\",2):f(\\\"\\\"{b=-i1nu@yp|ebUa7bM;gyt+:/ShNsozwzKtr2XaI5ub91+xzbt2M+6pTp<adbabQaHwD-jbP;QaDaz=8/db>yo7,bub0bB+r|\\\"\\\",2):f(\\\"\\\"}blbRycb,b0;p4y*Q/\\\"\\\",2):f(\\\"\\\"{|Jr0bbb:pH;rmX-g23,GyD=A;d|Na9*qhlb7b:44\\\"\\\",2):f(\\\"\\\"{kb\\\"\\\",2):f(\\\"\\\"{\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"{bdoc>\\\"\\\",2):f(\\\"\\\"}sw\\\"\\\",2):f(\\\"\\\"}7b\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}b1bEaTa|bvb-<w*8|\\\"\\\",2):f(\\\"\\\"{biqgnZ0v3Y;t3W;\\\"\\\",2):f(\\\"\\\"{bG2g9\\\"\\\",2):f(\\\"\\\"{bAak-Gy4iw*5,t20b<,3b;|7*56F,mb\\\"\\\",2):f(\\\"\\\"}+|b@aXaibRa4botizd|1bWatbcbVn=jn;Pa5+FaAaNaApOa136wSh-6rhp=@aRaS;6bjbttDaUa\\\"\\\",2):f(\\\"\\\"}=|20bE|2"));
$write("%s",("bfbH;ivfh?tt<*p@*Dtd</bNkPa+btqw\\\"\\\",2):f(\\\"\\\"{Mr2pQaxbU*8b/zA2fh3bB-T,nu?tMrs5<aUad:cbdbZaXqF+*b9b6pkbAalpebOaO*NgWa09lbd<UvDaTw=aG;ibJw+\\\"\\\",2):f(\\\"\\\"{9bkbTwubPa\\\"\\\",2):f(\\\"\\\"}/80-yd5tbrogbw1jb=afb/bt,cbz/yb@aO*|ikb=atle\\\"\\\",2):f(\\\"\\\"{2i1\\\"\\\",2):f(\\\"\\\"}0b<akb/7\\\"\\\",2):f(\\\"\\\"{be\\\"\\\",2):f(\\\"\\\"{4btqNaNgD\\\"\\\",2):f(\\\"\\\"}=.Y0=\\\"\\\",2):f(\\\"\\\"}o,M9xxyg=\\\"\\\",2):f(\\\"\\\"{-b<zwbVa9bzb=43b8r\\\"\\\",2):f(\\\"\\\"{bH1?a\\\"\\\",2):f(\\\"\\\"{b-1ubM+tb2zabV|njqw\\\"\\\",2):f(\\\"\\\"}wYyu811@aTa3yDxab?ybuib=a=j|8ibCu0b,bN|F44q5tubYaSwHsBam5k7jxajO|c,q9vb0\\\"\\\",2):f(\\\"\\\"{h|?3c\\\"\\\",2):f(\\\"\\\"{PaH+n-@tD9,ddb4b2\\\"\\\",2):f(\\\"\\\"{/zhbfb8ba|W-Jq,bQaCa@7wbP3MwSaOr5iVaM+@aybtb/08bJyAaytOahxPxFaSaYa\\\"\\\",2):f(\\\"\\\"{foyD+H9xx8bEa/9M+Za028ribh:jbB6=aWaPaI-hx>ajkc:a:2b:wzbu*f**bJp,\\\"\\\",2):f(\\\"\\\"}2.u2p2zb4bn*=avy"));
$write("%s",("RaJykb4w*bbbPtmbc4ub-lU0q,-l?.D\\\"\\\",2):f(\\\"\\\"}a1,5cjShY7>/.h=jOqgbmbFnA37bp3-b\\\"\\\",2):f(\\\"\\\"}xtwv-99,ia63b4|v8eb@7xu|bkx/bRaoweb*b7bOpQa4b,.cbI|u*aucbtb28=rdzP2jblbuv6b6pU-;u;7BnFa03*,cbTa|3\\\"\\\",2):f(\\\"\\\"}i.zrpk\\\"\\\",2):f(\\\"\\\"}6qbbybovdcJrVa8oCuXau|P7:wPaabxbQaZaU*TaKwbbbud0>a.b>aj-/bu/kbr28b51Op/bq+WaK+Fau\\\"\\\",2):f(\\\"\\\"}Bz4oV\\\"\\\",2):f(\\\"\\\"}<rE+y8|bRaBa\\\"\\\",2):f(\\\"\\\"{b1wYy*bStDwYaPr\\\"\\\",2):f(\\\"\\\"}xZaGx*bXaShk/Bwp5soWaN4*bJzX7mx+b8|8b8bq-IntbtbSatbWalb8b.+cbxb2tFa40hql\\\"\\\",2):f(\\\"\\\"{i\\\"\\\",2):f(\\\"\\\"{B7+57xu3ndmbhbj\\\"\\\",2):f(\\\"\\\"}3b+sDz2bBao|l-*0Bv4b4\\\"\\\",2):f(\\\"\\\"{th:,7,5b3bO|f7YadbP/81hbjb>a0bp7Da0b2bR|Ba2b9bZa9\\\"\\\",2):f(\\\"\\\"}3/k\\\"\\\",2):f(\\\"\\\"}?aCaTihbO|2b5bYadlFaCaLfNajbAaib/bhq4q-bBs+b5,F6r6q6vb2pm5a6UambH\\\"\\\",2):f(\\\"\\\"{g6mzAaI,Wa2..bxoEa\\\"\\\",2):f(\\\"\\\"}6A"));
$write("%s",("a=|2pVaTmSh=yEa<t|rVaRaEz/bSaQat2VarqO||b2b.bv2a|TaPr@aSa8b;hUag6WaRa?amb\\\"\\\",2):f(\\\"\\\"}0EaSambUaAaSaVaTaj+*bpolbubrykb2qcbAaL\\\"\\\",2):f(\\\"\\\"}:ou*6q?3ib>kgbD-@-FrTawbB*8h4bsp<5Fq;xbb6buhyb9b\\\"\\\",2):f(\\\"\\\"{wgpfbu,UuW4cbd1jkl\\\"\\\",2):f(\\\"\\\"{Iu\\\"\\\",2):f(\\\"\\\"}5>.Pur3abTtEwDq:1.rebpp|2+b@,Qs\\\"\\\",2):f(\\\"\\\"{bUaPa7b9zHzyby\\\"\\\",2):f(\\\"\\\"}y-fu0zk-ub3bE/:xSaabmb=a5bcb?akxryYapyu,Xap3Aamb+b.rWg3sCa<*7bb3Z201RtPtNtRamb|qdbQaq+hrMnw*bu4b7-t*8bBz?a8b>|Ksqo/0n/\\\"\\\",2):f(\\\"\\\"}bWpP+Fo-rFy<zDa2p5bVayb-bd1X\\\"\\\",2):f(\\\"\\\"{Sh=lVa?aOa*bcdztd1Fa..-bFa-\\\"\\\",2):f(\\\"\\\"}Jp3bhbYfZuYalzgkXaJru+bjXaubmb/t-tgtdblbp1GoBtHowr/bbbywv2oqSa>anuybK\\\"\\\",2):f(\\\"\\\"{Inwbhbuxib@aY-7p*,8b91E+fbabM\\\"\\\",2):f(\\\"\\\"}c/u\\\"\\\",2):f(\\\"\\\"}gnD\\\"\\\",2):f(\\\"\\\"}B.X0j\\\"\\\",2):f(\\\"\\\"{n,T0Da/b\\\"\\\",2):f(\\\"\\\"}sBaxbB*ybTa"));
$write("%s",("H-TaDa?ySh=*;*\\\"\\\",2):f(\\\"\\\"}x+bnj5bSaSa3j+bnutb|bpzWaAuPaScTaN*@ajtzdOaPaOaTz6bkb+bjbxbib12xt2pUa?aFx\\\"\\\",2):f(\\\"\\\"}bauZa=\\\"\\\",2):f(\\\"\\\"{ib\\\"\\\",2):f(\\\"\\\"}bjbfb,bCaBaKxrs10Zai+D16b4bebtqEaEaAaWaUa@vWaVaLwub>at+qqVa<0Xa:080-btpI1hbgbAv,p8b1\\\"\\\",2):f(\\\"\\\"{gbtbf1Y*t1\\\"\\\",2):f(\\\"\\\"}b/0s\\\"\\\",2):f(\\\"\\\"}+oNaAyYfAr0bowdxjyTm.v2\\\"\\\",2):f(\\\"\\\"}ub-bu1y//0Savb>aYa2plb3b\\\"\\\",2):f(\\\"\\\"}bQ0Sap15b/bub=awbtqtovyOaJy>aAuRaf*.b@a\\\"\\\",2):f(\\\"\\\"}bgb6bRabbbbfcBaTl|\\\"\\\",2):f(\\\"\\\"}j0r+7bh-+-wrJ0kbw*l\\\"\\\",2):f(\\\"\\\"{E\\\"\\\",2):f(\\\"\\\"}V0Nup,B\\\"\\\",2):f(\\\"\\\"}@.@\\\"\\\",2):f(\\\"\\\"}<.r+Pa|b|okv:gOae,OzZaUa6b8b7bho00,bUawu\\\"\\\",2):f(\\\"\\\"{pArIoab5bRtMfabgbwb4bd|2bDaw|ybhb>a7b3bEaU\\\"\\\",2):f(\\\"\\\"{lbSaqo=zs*fchqQa|\\\"\\\",2):f(\\\"\\\"}:\\\"\\\",2):f(\\\"\\\"{c-q+dbFaE,Ea@aEpmbr|9\\\"\\\",2):f(\\\"\\\"{=jcbFoWp9bEaVa|b<"));
$write("%s",("pbtC/A/?/lb\\\"\\\",2):f(\\\"\\\"}odb?rjbmbOaIrAaY\\\"\\\",2):f(\\\"\\\"}9oXa0*EaCa5s<pTaGne.Va2tZadymz,|8bN\\\"\\\",2):f(\\\"\\\"{0bFa9b6bL\\\"\\\",2):f(\\\"\\\"}tq4bYaSa\\\"\\\",2):f(\\\"\\\"{b*b3*Goqh1\\\"\\\",2):f(\\\"\\\"{YaPtSan.Mf*o\\\"\\\",2):f(\\\"\\\"{bzbCaCp7bmpBu.tWal/>a\\\"\\\",2):f(\\\"\\\"{bg*2pDafxAafu,qy\\\"\\\",2):f(\\\"\\\"{:z3b5bhbPa.b7br|/pgbXaBaybWa6bNac-<a*b\\\"\\\",2):f(\\\"\\\"}bxbPa6zEa5b0+Ergnl\\\"\\\",2):f(\\\"\\\"{3xXrm,Kul\\\"\\\",2):f(\\\"\\\"{r,l,,r3bdbp\\\"\\\",2):f(\\\"\\\"{Ca7mab0\\\"\\\",2):f(\\\"\\\"}n-Wa=aSa.bRa-vQaUq@a3b2p5,Ep5b0b1bT,O*db\\\"\\\",2):f(\\\"\\\"{bSa\\\"\\\",2):f(\\\"\\\"}bPaf-fb+,Wamb6bbcShJt5r1ba-hb9bly0b|bub9bu+4b2-2b+b?,I|8hKqRtVavxUaUaibac\\\"\\\",2):f(\\\"\\\"}bj+3b+bIroz4bXndc,byuebcx\\\"\\\",2):f(\\\"\\\"}bvb?adba-PnX*q-sjKzld*,\\\"\\\",2):f(\\\"\\\"}k*o\\\"\\\",2):f(\\\"\\\"}rTaTaWaUj3gibCaUq6bUalbSc0bdb\\\"\\\",2):f(\\\"\\\"}kzm@aZaBavbvbpzubzb@p\\\"\\\",2):f(\\\""));
$write("%s",("\\\"{vRa1bicSa9w*bmb*xTt1r.bWa?rvb7bFaZxSaybzbEaWaab2pzb/bBafb9b*bkbQa9b.bCa.b*b2bTaNa@aVaebbbboxbebZtUaWa,bXacb2b7bMnlbXtz+dxq*WabbEu.l>\\\"\\\",2):f(\\\"\\\"}Eu5xii?\\\"\\\",2):f(\\\"\\\"}C\\\"\\\",2):f(\\\"\\\"}ZaAajkWpf\\\"\\\",2):f(\\\"\\\"{C|cqGz|b\\\"\\\",2):f(\\\"\\\"}btbOamqdbvbshnvIyXue\\\"\\\",2):f(\\\"\\\"}QambebgzOaBa2prjErzbmzcb0zlbPaZa/bmz<aNaNpVa2b0q4igbXtyyQaJq0qQa1\\\"\\\",2):f(\\\"\\\"}mbp*,babXytbm*ubBa4bibzb?aUt3bcbebljtbwbTaVaEaShbxlbkbNa7yL*J*H*nhNaBa*b,b@a*b*bjbOazb<aL*tz-bOa0b,k2p0blb-b3sMrks<axxibWab*Qazb2pabwbOteb7bwbwbOafbRawb-rfw\\\"\\\",2):f(\\\"\\\"}bZaCaaqPaOpkbwykby\\\"\\\",2):f(\\\"\\\"{mb2pgb8bBaab.btb*p8bAajbgb0bjk-b,\\\"\\\",2):f(\\\"\\\"}*\\\"\\\",2):f(\\\"\\\"}|\\\"\\\",2):f(\\\"\\\"}FaxbkbWa5b-bvb+ugblbgpjuwr?xlbQa\\\"\\\",2):f(\\\"\\\"}xTaqh6bYaabab.zwb6bv\\\"\\\",2):f(\\\"\\\"{Eum\\\"\\\",2):f(\\\"\\\"{A\\\"\\\",2):f(\\\"\\\"}k\\\"\\\",2):f(\\\"\\\""));
$write("%s",("{enOubpgiZol\\\"\\\",2):f(\\\"\\\"{DulbNaVah|Mw=a8zPt,iTabbHszy0bvbVabbZamb\\\"\\\",2):f(\\\"\\\"{b4bovBaTapoh\\\"\\\",2):f(\\\"\\\"}7b+|5bovXaeb4u=vd\\\"\\\",2):f(\\\"\\\"{?\\\"\\\",2):f(\\\"\\\"{db=a7bDaebWuej\\\"\\\",2):f(\\\"\\\"}bfx1byuOa1zPaXa|b8b=akbgbuf,bkbbbwb3bZa1w0bmbybNa?aFa*bBw1s=v6btbib>adbib-d2pb|mbtb*b+b,bjyNkOz-b7ribSaX\\\"\\\",2):f(\\\"\\\"{.bowUa\\\"\\\",2):f(\\\"\\\"{bQaUa2b*b/bdz\\\"\\\",2):f(\\\"\\\"{bcb=aFaX27bhb/b|b,z*z<sabUa5btbgbFaOaWa0q0w2pBi@aFabb/bguXa@a9vtbfxytyb7\\\"\\\",2):f(\\\"\\\"{lbWa>rJybo\\\"\\\",2):f(\\\"\\\"}bibXa8bBsCaHzOaubcbEaRaAa3bLtVq0bQqWa|bab1z/z-z+zabPazbkb?a4vxbNa4b@aIq4bNaKt@w4bIogn4aHuh\\\"\\\",2):f(\\\"\\\"{Ju4x6xwbUabbzb*bYuIy<oQzSz0uhqrptbNa>aRahq.bNpPq=sdbVa;okblbvz2pwb*b|bBaub,i\\\"\\\",2):f(\\\"\\\"{zDakbEv<a9bxbbbPaIoGqcb/bwbSa1bZa|bWaubuvQaiy4bhbYaZaxbAa.bDa9b0bAaabYaDwgbbbMkBpwbEy8bebtoAa@v6ylbHwmb"));
$write("%s",("Eahx4b<agxmv+bVaCySaGxVaYaoywb?aGvOaXaRakbhbibcbib\\\"\\\",2):f(\\\"\\\"{b2p@azbRa0bWp4iDaZa2bqo5b>a=a2p2bAatbbb=aOa>aOpAaTaebSa3bubmxkxfbdbBvVa8biqbbVaOa,b\\\"\\\",2):f(\\\"\\\"}bPt,b9blbAagkyqxu3bjkbbibiqdbUa5w/bpx+bKxZw\\\"\\\",2):f(\\\"\\\"{qGa-s=a=aabibEaXa0bRa<aFa|s7bXaPaUa9bjbNaEuTr2xUrEu,lRrzxxxub9oCaotCaeb8bvxttNa1bPaPt>aNabb?aSa4i?aibab\\\"\\\",2):f(\\\"\\\"}b3bYacb7vgbabbb2b1b2p+b6bUwIr2p|bIr5sRaXaNa\\\"\\\",2):f(\\\"\\\"}wxbXatbXagt8bmbCa1b*b5tbblbibjbwblbXa4e*b=aYaRaabybOa7bgb5bCaUtSaub<axbEa0bcbQaTaiv7b\\\"\\\",2):f(\\\"\\\"{bub+b9byb2k5b4btbabtbBaibebclYaFa,b?qRvdsVaxbhqzbBq3j4iMp\\\"\\\",2):f(\\\"\\\"{bErnuYagrZaXanv<rZa7b.bhqej*p6b.bAq?azbsrtb\\\"\\\",2):f(\\\"\\\"{b/bcb@tXaDq*bbveb/bmbNazblb0bXaqvkbabcb7bBagbrj1bfb\\\"\\\",2):f(\\\"\\\"}b0b6p.b2tab4bgp=a-b/bfbQa|b/bUacbOa\\\"\\\",2):f(\\\"\\\"}bVq\\\"\\\",2):f(\\\"\\\"}b6gb"));
$write("%s",("b,rCagbCtPaeb>avbXaDa|bDa1bEucnLuGuZmapVrEuasWrYrhnZrQr3bFaybeb5bEaOs,sGa*s+udb3bPa6pDaRaybgbkbmbos<a<aub,rOaabtleb1bcbjbjkabep5bso,pyb7bZa>tfbcb0bfukbcbab2b8b0bZazb3jIttbSh?o8b/bXa>aub7btbdb*bEa2pSaUa|bkb2p9bvb,bRa7bNa.blbbbTaOoYa3b0q\\\"\\\",2):f(\\\"\\\"}bOaYa2k3bTacbGocbfbUa|ooq3jRa5bNaybfbfb1bubNa\\\"\\\",2):f(\\\"\\\"}bVatbfbwbebhbwsxb8bFaibib4b2pyblbTagbZbjbRaWaLpFa\\\"\\\",2):f(\\\"\\\"}bzb7b5swbCa2pibQq8b.b8oPrcb|i2pYaeb.b=a4bKoFa\\\"\\\",2):f(\\\"\\\"{s-bbbuqybbrxbMf|q5bOa3bQa7bRaCaShgsJqShHq@a/bPaPa*bmoUagq=r3jVaUaTaBacbmbrofbvb0b0b2p-bXakbCaDigngiXoSrYocpWogngn;iQoXambzb@a-bfb|b6b,b3jmbjbcb,rIo8babXaablb\\\"\\\",2):f(\\\"\\\"{b-bzbMf>aebvbTa1b3j\\\"\\\",2):f(\\\"\\\"{b1bkb9b\\\"\\\",2):f(\\\"\\\"{rebzbNaubQa\\\"\\\",2):f(\\\"\\\"{b.b?aab@pabFaRa\\\"\\\",2):f(\\\"\\\"}bTaYa-bWa+bBaTg4eKqIqGqVa-bwbBqQaybDa@aSh1p\\\"\\\""));
$write("%s",(",2):f(\\\"\\\"{bebYaQa8b\\\"\\\",2):f(\\\"\\\"{f>a+b2q6b-b9bfb-b3bUa2p7bVaXa5b7b2b0bPayqwq*bNahbUavb@aGpvbZaaqmb|odbub\\\"\\\",2):f(\\\"\\\"}bkbdbmb4bTa<a7bdb0bKoWaxb2p,blbUaQa>a|oebVajbjb7b0bWaBaFa+bSawb@aUa5peb:pqpsoBaDazb=aEihb*bBambPa0bEajbFaPaCambFa>aTafbibOaCajbhb6bXaHo3b7p+dXabb\\\"\\\",2):f(\\\"\\\"}bxgGa@oPa4bvbcbwb=a,bZahbslcb@atb>aLojbtckbibDaFa5b1bDawb5b\\\"\\\",2):f(\\\"\\\"}bCa4bso0bibvbiiSoTo|lRo|lUofniijnkniiingnxo-b6fjbPa,btkwbmbSaXaFa6b/b\\\"\\\",2):f(\\\"\\\"}bShqbAa-bCaFa-b7bTaQaRnYaaomb,bYa-o.o,o*o7b/bYagbib,bjbvbRaQa|diboi|bmbXaZa\\\"\\\",2):f(\\\"\\\"{b?enkEahoTaRa>aFasgybdb.b3jeblbzb,bNa7bvbCaEahb<aCabb*bWgQaub*bWaQagbSa,bEa7b6bAaEaHl7nvn;mkmimonEfQmsmqm-n;a>mrmpmQm=m:l\\\"\\\",2):f(\\\"\\\"{n-bHl4mCa9lNmwbicQm;lhmrnEaSl>mjm9lxmemcmgn0l0lan4adn9agibn|lYm+lii/l/b\\\"\\\",2):f(\\\"\\\"{f-a|hub.h8a5mB"));
$write("%s",("mymGm8l9aEaOa>m<m-m8f:a-b>m=aAa-a.m|mCaSlWlwm@a<a-b|e1m\\\"\\\",2):f(\\\"\\\"{mKlgmVlMlKlIlnmzm:aCa|etm>aAahmRlMl9a6lNlAa?a>aDl|efmslHlUlBa-aJlClAl*bvbtb/b-a+bId<lOl=lFl@aDlHlSe|eBlGl?aAa9l\\\"\\\",2):f(\\\"\\\"{b7l>l<lFa:l8l6lHa4l9a|e5lxb8a+e-a1bLf8aEfpl8arb|eidfi-l-l\\\"\\\",2):f(\\\"\\\"}l3a:igi\\\"\\\",2):f(\\\"\\\"{l-fhiil<h7f6b-a+czbxbubHaqb6aqb3i4i2i5aqb-g-aff1bzb.b6fnbxbkiShHgFghgHfkhxhbkxjZj?a=a:i;d\\\"\\\",2):f(\\\"\\\"}h2kyiIjdh.ktcBa3a=h6g2iwb=fTjakFjBa?a9i6e|hrbLj?aJjSjviGjDa?aDj2b3b5iBf+c:g-a8f-b1jCa3aKa\\\"\\\",2):f(\\\"\\\"{b;atgwbccIa3b1bnj,b|b0adhyhdhzjRjvjCa9i.bbi?a?iyj=i;i@a9iyb3bBjyh2h>iwhwjBa>a9iPcsihghgsbubwbSh-a2j0j:a;b-j1b0b-b3aAa3a7b-aSh.a:b:b,byhlhxiPaUh<i@a3a|hwb+b-aPcbj/b8b1bPcxb;aBf-b;gZaWf|b.b5b-aTi,i3bDfvb|b6g5iWfMf3bgf;a<b:b3b-a8b6g,bxb2b2btb;ayhEhwiEh3a>a3a5anb-a3i/b3b"));
$write("%s",("4b.bHa8byb2bsgtbDfxb5b+bGgyhwhThGhlh?g8f6fHaoioiFaGaRh|fld4aogei/ach4a-aMfKfMaFa=aEh-bGh2h1hGa+bJd?h9a/b5a|fCcyg-bPaBaob2h6aKaMa9aMaIa5axb3b.b4b0bxb*htbLfyhRfwhGaMb5g2bzb;azb-b7fccJaWg?achlhCdYaOaVafbVaibNa=adhdh?a;aAgVaNaUaogchRfvbpbEa*c7b?aDaBaCa>anbJdubSczb=fIc?gyfwfuf2bsfNd3bHa?e-a-fGf:aIa+ctb,b:avbldub4bcb-btggcqgHaebdbJaGagfef8a1bxbwbtbxbUaac|b3bKffb/aRfggtbxc?f?a1aRf-a6a5bOf>azd:a,cNaOfwb.b;b>aHfob,c:a-a.b\\\"\\\",2):f(\\\"\\\"{bvbxb5a1aob,fCe2b-a:b1dtbHa6a/c2b/a:f-f;d+c1b/b3dMd-aDdBd@dmf/aob5a.d,d*d-b4b7eSc;axb+b.bbcZb0cbfJasdHa/aed+e0cGb/d,btb-b4aWbudpcgdLc=chchd6areOapc0cNb/a;bje/eGaHb5dedOb.a8aNd8aLdLa=a>aIaOaJapb6a+e5azb+cdcfbhc;aOaFdYd6aHaCa@aIaQd8aHa=a.cIbCbMd\\\"\\\",2):f(\\\"\\\"{cycvcocRapcXbocTa;b;bpbgbYdJaGbRanbQaJagbnbcb>dqc5dpbebnbOa8a0c4aJaTa5a+btb5"));
$write("%s",("bxbJaQa,c*cRa5a1bzc6aedMa0c3bldjd;aeded8ard5a6a5aedxb/btbvb2bxb,c1b4b3bxb1b0cocPa8aNapcMagdUc3b|b+b/b2b4arcFbnc4a=a?axbtc4aSbJcPbKckcic+bZb3b-bzcXbqcFb5aMa/ancvc+b+b|byb4a9cVbNa5aRb7cFbnbFbMapb2c.aMaFb.a4a5aJaOa-a-b|b-aeb5aicybHa<b/akc>a>aXb6aOb/a8a6a/apb4a1b.b3bvb4b1b3b2b-b.bvb4anb/aJaPa5a8a4a6apbEb5a5aBb,b9a4apbpbnb8anb4aGa=a:bJacb!\\\"\\\",2):f(\\\"\\\"})23(f\\\"\\\",2):f(\\\"\\\"{#~[2xha=s,y=z,13&X3^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'yay,]99999[gnirtS wen=][c n3aea\\\"\\\",2):f(\\\"\\\"{)v]y3b&a(niam diov citats cilbup\\\"\\\",2):f(\\\"\\\"{RQ ssalcz4rfa cdlnl3c/a;maertStnirP/oi/avajL tuo/metsyS/gn"));
$write("%s",("al/avajm4bdateg@3doa2 kcats timil.v3dga]; V);Q4aC3ecaL[b5aX4hha dohtem?3e;4nga repus&3ecaRQ@3cgassalc.<5joa(=:s;0=:c=:i;)|4ajaerudecorp/3f\\\\\\\"\\\"),\\\\n(\\\\\\\"\\\"qa(tnirp.biL.oken\\\"\\\",2):f(\\\"\\\"{.3bianoitcnufR6\\\"\\\",2):f(\\\"\\\"{sa(rtStup=niam^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^127^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^32^[2fha\\\"\\\",2):f(\\\"\\\"})1(f\\\"\\\",2):f(\\\"\\\"{#v3mja51(f\\\"\\\",2):f(\\\"\\\"{#,4353(ga13(f\\\"\\\",2):f(\\\"\\\"{#j4[j4boa(etirw.z;)tuo.N8aba(67b~auptuOPIZG.piz.litu.avaj wen=zG4Zka30341(f\\\"\\\",2):f(\\\"\\\"{#tm4[m4c5aR0Z0Z/512152353/2/2166263="));
$write("%s",("4/3141726??:1518191:1/@4[@4cda*6 Q5[p4dea1312^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'5[w8[$5ofa41310r4[r4c7=[B>[j4[^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'6pma(amirpmi oicy4[(5[j4hma++]371[]591[?6[?6cpani;RQ omtirogla\\\"\\\",2):f(\\\"\\\"{4[\\\"\\\",2):f(\\\"\\\"{4cCa;t:\\\"\\\",2):f(\\\"\\\"}%%%%\\\"\\\",2):f(\\\"\\\"}fi\\\"\\\",2):f(\\\"\\\"}*-84\\\"\\\",2):f(\\\"\\\"})48361(f\\\"\\\",2):f(\\\"\\\"{#]i[\\\"\\\",2):f(\\\"\\\"{\\\"\\\",2):f(\\\"\\\"}+17\\\"\\\",2):f(\\"));
$write("%s",("\"\\\"{<84.;i:-i602\\\"\\\",2):f(\\\"\\\"{;i:911\\\"\\\",2):f(\\\"\\\"{;j:632*7[ra116(f\\\"\\\",2):f(\\\"\\\"{#(tnirP.tmfIIcfacnuf;&4[&4bdatmfn4[n4cgaropmi;ILagagakcap~4Zea5102T6dbapD6[r4cba-l4[l4bpatnirp tesn\\\"\\\",2):f(\\\"\\\"})420aEaka etalpmet.r8[ma99(f\\\"\\\",2):f(\\\"\\\"{#(ntnire8[ia974(f\\\"\\\",2):f(\\\"\\\"{#fp4[ga^64^\\\"\\\",2):f(\\\"\\\"})32u9awa,s(llAetirW;)(resUtxeTOPada=:s%8[ba9#8eo4[ia9(f\\\"\\\",2):f(\\\"\\\"{#S Cm4[-Eaca&(y5[ga9(f\\\"\\\",2):f(\\\"\\\"{# .6[.6[.6oiaRQ margo&5[t4cjaS D : ; R-5[6L[j4[j4o%6[k4aqa. EPYT B C : ; Az4[56[j4[j4nka)*,*(ETIRW/6[J7chaA B : ;s4[s4aba [2cr4[*5dia: ^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"' "));
$write("%s",("ohce3B[EYaeastupLRcdatniy4/ca0153.ea%%%%m4[m4[53ipaparwyyon noitpoz4023[230ca(nRO.%a7(f\\\"\\\",2):f(\\\"\\\"{#(etirwf:oin\\\"\\\",2):f(\\\"\\\"})4(f\\\"\\\",2):f(\\\"\\\"{#>-)_(niamp3cvP)ka(f\\\"\\\",2):f(\\\"\\\"{# cnirp,L)k;eja.OI[p]^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'[(3rba@2Wa6;alaM dohtem06x*3c|5aU;cpadiov;oidts.dts 6Yab4kkaenil-etirwb5dva(,^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\""));
$write("%s",("\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'s%^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'(gol.elosnoc;)^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'73g\\\"\\\",2):f(\\\"\\\"}a^129^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f"));
$write("%s",("(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"' nioj.)1+n(yarrA>-)n(=fI3cwa^31^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",2):f(\\\"\\\"}54,1\\\"\\\",2):f(\\\"\\\"{.^127^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"# qes-er()|3cH3bba^31^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"p3lg3fw3hla1% ecalper.j4dea^128^jAc/arts(# pam(]YALPSID^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^127^\\\"\\\",57):"));
$write("%s",("f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\".NOISIVID ERUDECORPA3cma.RQ .DI-MARGv3g53d|bNOITACIFITNEDI^127^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"[tac-yzal(s[qesod(^63^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"))System.Console.Write($^63^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"Put caffeine \\\"\\\",2):f(\\\"\\\"{(int)c\\\"\\\",2):f(\\\"\\\"} into the mixing bowl.^64^n^63^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\");M3pva^63^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"Liquify contents ofE3oeaPour^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):"));
$write("%s",("f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'3w^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^1^\\\"\\\",4):f(\\\"\\\"'4e\\\"\\\",2):f(\\\"\\\"{abaking dish.^64^n^64^nServes 164cma\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}^31^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\");\\\"\\\",2):f(\\\"\\\"}/****/e3a^15^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"),s[999999],*q=s;int main()\\\"\\\",2):f(\\\"\\\"{int n,m;for(;*p;)\\\"\\\",2):f(\\\"\\\"{n=(*p-5)%9"));
$write("%s",("2+(p[1]-5)%92*87;p+=2;if(n>3999)for(m=(*p++-5)%92+6;m--;q++)*q=q[4000-n];else for(;n--;)*q++=*p++;\\\"\\\",2):f(\\\"\\\"}puts(s);return 0;\\\"\\\",2):f(\\\"\\\"}^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"))\\\"\\\",2):f(\\\"\\\"{s+=^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"00g,^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\";for(m=1;m<256;m*=2)s+=^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"00g,4,:^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"+(c/m%2>0?^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"4+^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\""));
$write("%s",("\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\":^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\")+^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\",^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\";f(s);s=^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"4,:,^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\";\\\"\\\",2):f(\\\"\\\"}f(s+s);for(c:Base64.getDecoder().decode(^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"kaAREREX/I0ALn3n5ef6l/Pz8+fnz58/BOf5/7/hEX/OZzM5mCX/OczmZ"));
$write("%s",("zBPn5+X/OczMznBL/nM5mZzBPu++fPPOc5zngnnOZzOZgnBMGAW7A==^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"))\\\"\\\",2):f(\\\"\\\"{c=c<0?256+c:c;for(i=0;i++<3;c/=8)f(c%8);f(^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"8*+8*+,^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\");\\\"\\\",2):f(\\\"\\\"}f(^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"@^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\");^1^\\\"\\\",4):f(\\\"\\\"'|sed -e^1^\\\"\\\",4):f(\\\"\\\"'s/^16^/^32^/g^1^\\\"\\\",4):f(\\\"\\\"' -e^1^\\\"\\\",4):f(\\\"\\\"'s/^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"/^16^q/g^1^\\\"\\\""));
$write("%s",(",4):f(\\\"\\\"' -e^1^\\\"\\\",4):f(\\\"\\\"'s/.*/print ^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&^7^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"^8^nquit/^1^\\\"\\\",4):f(\\\"\\\"'^3^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\")\\\"\\\",2):f(\\\"\\\"}^1^\\\"\\\",57):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\")\\\"\\\",4):f(\\\"\\\"');\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\").split(\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",64):f(\\\"\\\"^\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\");for(int i=1;i<a.length;a[0]+=a[i+1],i+=2)\\\"\\\",2)"));
$write("%s",(":f(\\\"\\\"{a[0]+=\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",89):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\".repeat(Integer.parseInt(a[i]));\\\"\\\",2):f(\\\"\\\"}System.out.print(a[0]);\\\"\\\",2):f(\\\"\\\"}\\\"\\\",2):f(\\\"\\\"}\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\";FORiTO UPBtDO INTn:=ABSt[i];print(REPR(50+n%64)+c+REPR(50+n%8MOD8)+c+REPR(50+nMOD8)+b+\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"J\\\"\\\",25):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"+a)OD\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\")\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"while(!=(S:length)0)\\\"\\\",2):f(\\\"\\\"{\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"trans c(S:read)\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\""));
$write("%s",(",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"D(c:to-integer)\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"f 35 39\\\"\\\",2):f(\\\"\\\"}\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"f 24 149\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"interp:library\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"afnix-sio\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"trans o(afnix:sio:OutputTerm)\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"&Character\\\"\\\",4):f(\\\"\\\"'Val(10)&\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\"o:write B\\\"\\\",9):f(\\\"\\\"\\\\\\\"\\\");end;\\\"\\\",1):f(\\\"\\\"\\\\\\\"\\\")\\\"\\\",1):f(\\\"\\\"nsys.exit 0'}\\\\\\\"\\\")\\\"\\\",0)]]></xsl:template></xsl:stylesheet>\\\":s=\\\"   \\\":For i=0To 7:s &=Chr(32-(Asc(c)>>7-i And"));
$write("%s",(" 1)*23):Next:System.Console.Write(s &n &Chr(9)&n &\\\"  \\\"):Next:System.Console.Write(n &n &n):End Sub:End Module\")\nput=s\nprint\nqa!"));
end endmodule